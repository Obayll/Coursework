--------------------------------------------------------------------------------------------
-- Course: ECE 332 - Digital System Design Lab
-- Author: 
-- 
-- Create Date: 
-- Experiment Name: Arithmetic and Logic Unit in VHDL (Lab #8)
-- Project Name: project_8 - Behavioral
--
-- Description:	Test bench for the 4-bit Arithmetic and Logic Unit.
-- 				It tests all 12 ALU operations.
--				For the binary operations, it tests four combinations of the inputs: +/+, +/-, -/+, and -/-
--				For the unary operations, it tests a + input and a - input.
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
-- Insert additional package here (if needed).

entity project_8_tb is
end project_8_tb;

architecture behavior of project_8_tb is

-- Insert component declaration for device under test (DUT) here.

-- Insert signal declarations here.

begin

-- Insert component instantiation (i.e. port map statement) here.
	
	ALU_simulation : process
	begin

	-- Insert your testbench code here.

	end process ALU_simulation;
	
end behavior;
