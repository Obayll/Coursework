--------------------------------------------------------------------------------------------
-- Course: ECE 332 - Digital System Design Lab
-- Author: 
-- 
-- Create Date: 
-- Experiment Name: Arithmetic Circuits in VHDL (Lab #6)
-- Project Name: project_6 - Behavioral
--
-- Description:	Test bench for the 4-bit Adder in Project_6 (Lab_6_2).
--				It tests all 2^4 x 2^4 = 256 combinations of the inputs.
--				This is known as an "exhaustive test".
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
-- Insert additional package here.

entity project_6_tb is
end project_6_tb;

architecture behavior of project_6_tb is

-- Insert component declaration for device under test (DUT) here.

-- Insert signal declarations here.

begin

-- Insert component instantiation (i.e. port map statement) here.
	
	Adder_simulation : process
	begin

	-- Insert your testbench code here.
	
	end process Adder_simulation;
	
end behavior;
